`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/08/07 15:54:12
// Design Name: 
// Module Name: Asyfifo_data_stream_ctr
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Asyfifo_data_stream_ctr
#(parameter DATA_SIZE  = 16 ,//data width                                                                
  parameter DEPTH_SIZE = 10 ,//data depth 2^DEPTH_SIZE(10:1024)                                          
  parameter FULL_THR   = 512,//user define full threshold assert value                                   
  parameter FULL_THR_EN= 1  ,//0/1:disable/enable user define full threshold assert value                
  parameter WR_CLK_PR  = 20 ,                                                                              
  parameter RD_CLK_PR  = 8                                                                                
)
(   //input sign
    input                       rst_n          ,
    //push data in ctr
    input                       clk_in         ,
    input     [DATA_SIZE-1:0]   data_in        ,
    input                       data_in_en     , 
    //pop data out ctr         
    input                       clk_out        ,
    input                       data_out_en    ,//data out requst
    //output sign
    output reg                  data_out_ready ,//any fifoN had full or prog_full   
    output reg                  data_out_busy  ,  
    output reg [DATA_SIZE-1:0]  data_out       
    );
 
//localparam  DATA_DEPTH = 1024;    
localparam  DATA_DEPTH =  2**DEPTH_SIZE;  

//fifo1 and fifo2 port define
wire                  data1_in_en   ; 
wire                  data2_in_en   ;    
wire                  data1_out_en  ; 
wire                  data2_out_en  ; 
wire [DATA_SIZE-1:0]  data1_out     ;
wire [DATA_SIZE-1:0]  data2_out     ; 
wire                  fifo1_full    ;
wire                  fifo2_full    ;  
wire                  fifo1_empty   ;
wire                  fifo2_empty   ;
wire [DEPTH_SIZE:0]   rd_data1_count;  
wire [DEPTH_SIZE:0]   rd_data2_count;
wire [DEPTH_SIZE:0]   wr_data1_count;
wire [DEPTH_SIZE:0]   wr_data2_count;   
wire                  prog1_full    ;
wire                  prog2_full    ;


//data push into fifo 
localparam st_push_idle        = 5'b00001;
localparam st_push_fifo1       = 5'b00010;
localparam st_push_fifo2_wait  = 5'b00100;//wait fifo2 had pop
localparam st_push_fifo2       = 5'b01000;
localparam st_push_fifo1_wait  = 5'b10000;//wait fifo1 had pop

reg [4:0] cur_push_state;
reg [4:0] nex_push_state;


//data pop from fifo
localparam st_pop_idle   = 3'b001;
localparam st_pop_fifo1  = 3'b010;
localparam st_pop_fifo2  = 3'b100;
reg [2:0] cur_pop_state;
reg [2:0] nex_pop_state;
//data in fifo en
assign data1_in_en = (cur_push_state == st_push_fifo1)?data_in_en:1'b0;
assign data2_in_en = (cur_push_state == st_push_fifo2)?data_in_en:1'b0;
//data out fifo en
assign data1_out_en = (cur_pop_state==st_pop_fifo1)?data_out_en:1'b0;
assign data2_out_en = (cur_pop_state==st_pop_fifo2)?data_out_en:1'b0;

always@(*)begin
    if(!rst_n)begin
        data_out = {DATA_SIZE{1'b0}};
    end
    else if(data_out_busy)begin
        if(cur_pop_state==st_pop_fifo1)begin
            data_out = data1_out;
        end
        else if(cur_pop_state==st_pop_fifo2)begin
            data_out = data2_out;
        end
        else begin
            data_out = data_out;
        end  
    end  
    else begin
        data_out = {DATA_SIZE{1'b0}};
    end
end

//assign data_out = (((cur_pop_state == st_pop_fifo1)||(cur_pop_state == st_pop_fifo2))&&(data_out_busy))? ((cur_pop_state == st_pop_fifo1)? data1_out:data2_out):{DATA_SIZE{1'b0}};
//assign data_out = (((cur_pop_state == st_pop_fifo1)||(cur_pop_state == st_pop_fifo2)))? ((cur_pop_state == st_pop_fifo1)? data1_out:data2_out):{DATA_SIZE{1'b0}};
//data push into fifo(State transitions) 
always@(posedge clk_in or negedge rst_n)begin
    if(!rst_n)begin
        cur_push_state <= st_push_idle  ;    
    end
    else begin
       cur_push_state  <= nex_push_state;  
    end
end



always@(*)begin
    nex_push_state <=  st_push_idle;
    case(cur_push_state)
        st_push_idle:begin
                nex_push_state <= st_push_fifo1;
        end
        st_push_fifo1:begin
            if((FULL_THR_EN&&prog1_full)|fifo1_full)begin
                if(fifo2_empty)
                    nex_push_state <= st_push_fifo2;
                else
                    nex_push_state <= st_push_fifo2_wait;
            end    
            else begin
                nex_push_state <= st_push_fifo1;         
            end
        end    
        st_push_fifo2_wait:begin
            if(fifo2_empty)begin
                nex_push_state <= st_push_fifo2;           
            end    
            else begin
                nex_push_state <= st_push_fifo2_wait;
            end
        end 
        st_push_fifo2:begin
            if((FULL_THR_EN&&prog2_full)|fifo2_full)begin
                if(fifo1_empty)
                    nex_push_state <= st_push_fifo1;
                else
                    nex_push_state <= st_push_fifo1_wait;
            end    
            else begin
                nex_push_state <= st_push_fifo2;         
            end
        end    
        st_push_fifo1_wait:begin
            if(fifo1_empty)begin          
                nex_push_state <= st_push_fifo1;
            end    
            else begin
                nex_push_state <= st_push_fifo1_wait;
            end
        end
        default:begin
            nex_push_state <= st_push_idle;
        end         
    endcase
end

//data pop into fifo(State transitions) 
always@(posedge clk_out or negedge rst_n)begin
    if(!rst_n)begin
        cur_pop_state  <= st_pop_idle  ;    
    end
    else begin
        cur_pop_state  <= nex_pop_state;  
    end
end


always@(*)begin
    nex_pop_state <= st_pop_idle;    
    case(cur_pop_state)
        st_pop_idle:begin
            if(prog1_full|fifo1_full)begin          
                nex_pop_state <= st_pop_fifo1;
            end
            else if(prog2_full|fifo2_full)begin        
                nex_pop_state <= st_pop_fifo2;
            end    
            else
                nex_pop_state <= st_pop_idle;     
        end
        st_pop_fifo1:begin
            if(!fifo1_empty)begin
                nex_pop_state <= st_pop_fifo1;
            end    
            else begin
                nex_pop_state <= st_pop_idle;
            end
        end  
        st_pop_fifo2:begin
            if(!fifo2_empty)begin
                nex_pop_state <= st_pop_fifo2;
            end    
            else begin
                nex_pop_state <= st_pop_idle;
            end
        end 
        default:begin
            nex_pop_state <= st_pop_idle;
        end 
    endcase
end

always@(posedge clk_out or negedge rst_n)begin
    if(!rst_n)
        data_out_ready <= 1'b0;
    else if(((wr_data1_count==FULL_THR)&prog1_full)|((wr_data2_count==FULL_THR)&prog2_full)
            |((wr_data1_count==DATA_DEPTH)&fifo1_full)|((wr_data2_count==DATA_DEPTH)&fifo2_full))
        data_out_ready <= 1'b1;
    else    
        data_out_ready <= 1'b0;
end

//data_out_busy
reg data_out_busy_en;
always@(posedge clk_out or negedge rst_n)begin
    if(!rst_n)begin
        data_out_busy    <= 1'b0;
        data_out_busy_en <= 1'b0;
    end
    else begin
        if((cur_pop_state==st_pop_fifo1)|(cur_pop_state==st_pop_fifo2))begin
            if(data_out_en)begin
                data_out_busy_en <= 1'b1;
                //data_out_busy <= 1'b1;
            end
            if(data_out_busy_en)
                data_out_busy <= 1'b1;
        end
        else begin
            data_out_busy <= 1'b0;   
            data_out_busy_en <= 1'b0;
        end 
    end
end

async_fifo 
#(.DATA_SIZE  (DATA_SIZE  ),//data width
  .DEPTH_SIZE (DEPTH_SIZE ),//data depth 2^DEPTH_SIZE(10:1024)
  .FULL_THR   (FULL_THR   ),//user define full threshold assert value
  .FULL_THR_EN(FULL_THR_EN))//0/1:disable/enable user define full threshold assert value 
u0_async_fifo(
    //input sign  
     .rst_n        (rst_n         ),//input                ��λ
     .wr_clk       (clk_in        ),//input                дʱ�� 
     .wr_en        (data1_in_en   ),//input                д��ʹ��                      
     .din          (data_in       ),//input [DATA_SIZE-1:0]д������
     .rd_clk       (clk_out       ),//input                ��ʱ��                 
     .rd_en        (data1_out_en  ),//input                ����ʹ�� 
    //output sign
     .dout         (data1_out     ),//output [DATA_SIZE-1:0]��������
     .full         (fifo1_full    ),//output                д���ź�
     .empty        (fifo1_empty   ),//output                �����ź�   
     .rd_data_count(rd_data1_count),//output [DEPTH_SIZE:0] �ɶ�������        
     .wr_data_count(wr_data1_count),//output [DEPTH_SIZE:0] ��д������        
     .prog_full    (prog1_full    ) //output                �ﵽFULL_THR���ź�
    );    
    
async_fifo 
#(.DATA_SIZE  (DATA_SIZE  ),//data width
  .DEPTH_SIZE (DEPTH_SIZE ),//data depth 2^DEPTH_SIZE(10:1024)
  .FULL_THR   (FULL_THR   ),//user define full threshold assert value
  .FULL_THR_EN(FULL_THR_EN))//0/1:disable/enable user define full threshold assert value 
u1_async_fifo(
    //input sign  
     .rst_n        (rst_n         ),//input                ��λ
     .wr_clk       (clk_in        ),//input                дʱ�� 
     .wr_en        (data2_in_en   ),//input                д��ʹ��                      
     .din          (data_in       ),//input [DATA_SIZE-1:0]д������
     .rd_clk       (clk_out       ),//input                ��ʱ��                 
     .rd_en        (data2_out_en  ),//input                ����ʹ�� 
    //output sign
     .dout         (data2_out     ),//output [DATA_SIZE-1:0]��������
     .full         (fifo2_full    ),//output                д���ź�
     .empty        (fifo2_empty   ), //output                �����ź� 
     .rd_data_count(rd_data2_count),//output [DEPTH_SIZE:0] �ɶ�������        
     .wr_data_count(wr_data2_count),//output [DEPTH_SIZE:0] ��д������        
     .prog_full    (prog2_full    ) //output                �ﵽFULL_THR���ź�
    );     

    
endmodule
