`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/08/08 15:36:29
// Design Name: 
// Module Name: define
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define DATA_SIZE    16 
`define DEPTH_SIZE   10 
`define DATA_DEPTH   2**10
`define FULL_THR     512
`define FULL_THR_EN  1  
`define WR_CLK_PR    20                                                                             
`define RD_CLK_PR    8  
